module tb();

mipsprocessor hamada ();

endmodule 

// 
