module  adder (pc, newpc);

 
input [31:0] pc;

output[31:0] newpc;


wire [31:0] pc;

wire [31:0] newpc;


assign newpc=pc+4 ;

 
endmodule 
  
